library verilog;
use verilog.vl_types.all;
entity Proposed_Tb is
end Proposed_Tb;
